module halfadder(A,B,sum,c_out);

	input A,B;
	
	output sum,c_out;
	
	xor IC7486(sum,A,B);
	and IC7408(c_out,A,B);
	
endmodule